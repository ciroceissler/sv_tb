interface tb_if;
interface : tb_if
