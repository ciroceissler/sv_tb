class test_base;
endclass : test_base
