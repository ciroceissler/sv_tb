class test_rand2;
endclass : test_rand2
