class agent;
  function new();
  endfunction : new

  task run();
  endtask : run
endclass
