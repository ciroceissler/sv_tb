class packet;
  function new();
  endfunction : new
endclass
