class scoreboard;
  function new();
  endfunction : new
endclass
