module testbench;
endmodule : testbench
