class test_rand1;
endclass : test_rand1
