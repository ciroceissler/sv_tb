class monitor;
  function new();
  endfunction : new
endclass
