module dut();
endmodule : dut
