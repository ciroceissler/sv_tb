program run_test();
endprogram : run_test
